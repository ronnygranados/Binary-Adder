module adder(a, b, cin, q, cout);

    // Comments

endmodule